LIBRARY ieee;
USE ieee.std_logic_1164.ALL;

ARCHITECTURE behavior OF mips_processor  IS


